library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;


entity dram is
    generic ( maxAddrBit : integer := 8;
              wordSize   : integer := 16
            );
    port (clk             : in  std_logic;
          areset          : in  std_logic;
          mem_writeEnable : in  std_logic;
          mem_readEnable  : in  std_logic;
          mem_addr        : in  std_logic_vector(maxAddrBit-1 downto 0);
          mem_write       : in  std_logic_vector(wordSize-1 downto 0);
          mem_read        : out std_logic_vector(wordSize-1 downto 0);
          mem_busy        : out std_logic
        );
end dram;

architecture dram_arch of dram is


type ram_type is array(natural range 0 to (2**maxAddrBit)-1) of std_logic_vector(wordSize-1 downto 0);

shared variable ram : ram_type := (
0 => x"0000",
1 => x"0170",
2 => x"02e0",
3 => x"044f",
4 => x"05be",
5 => x"072c",
6 => x"0898",
7 => x"0a04",
8 => x"0b6e",
9 => x"0cd6",
10 => x"0e3c",
11 => x"0fa0",
12 => x"1102",
13 => x"1261",
14 => x"13bd",
15 => x"1516",
16 => x"166c",
17 => x"17be",
18 => x"190d",
19 => x"1a58",
20 => x"1b9e",
21 => x"1ce1",
22 => x"1e1f",
23 => x"1f58",
24 => x"208d",
25 => x"21bd",
26 => x"22e7",
27 => x"240c",
28 => x"252b",
29 => x"2645",
30 => x"2759",
31 => x"2867",
32 => x"296e",
33 => x"2a6f",
34 => x"2b6a",
35 => x"2c5e",
36 => x"2d4b",
37 => x"2e31",
38 => x"2f10",
39 => x"2fe7",
40 => x"30b8",
41 => x"3180",
42 => x"3241",
43 => x"32fb",
44 => x"33ac",
45 => x"3456",
46 => x"34f7",
47 => x"3591",
48 => x"3622",
49 => x"36aa",
50 => x"372b",
51 => x"37a2",
52 => x"3812",
53 => x"3878",
54 => x"38d6",
55 => x"392b",
56 => x"3977",
57 => x"39bb",
58 => x"39f5",
59 => x"3a27",
60 => x"3a4f",
61 => x"3a6f",
62 => x"3a85",
63 => x"3a93",
64 => x"3a97",
65 => x"3a93",
66 => x"3a85",
67 => x"3a6f",
68 => x"3a4f",
69 => x"3a27",
70 => x"39f5",
71 => x"39bb",
72 => x"3977",
73 => x"392b",
74 => x"38d6",
75 => x"3878",
76 => x"3812",
77 => x"37a2",
78 => x"372b",
79 => x"36aa",
80 => x"3622",
81 => x"3591",
82 => x"34f7",
83 => x"3456",
84 => x"33ac",
85 => x"32fb",
86 => x"3241",
87 => x"3180",
88 => x"30b8",
89 => x"2fe7",
90 => x"2f10",
91 => x"2e31",
92 => x"2d4b",
93 => x"2c5e",
94 => x"2b6a",
95 => x"2a6f",
96 => x"296e",
97 => x"2867",
98 => x"2759",
99 => x"2645",
100 => x"252b",
101 => x"240c",
102 => x"22e7",
103 => x"21bd",
104 => x"208d",
105 => x"1f58",
106 => x"1e1f",
107 => x"1ce1",
108 => x"1b9e",
109 => x"1a58",
110 => x"190d",
111 => x"17be",
112 => x"166c",
113 => x"1516",
114 => x"13bd",
115 => x"1261",
116 => x"1102",
117 => x"0fa0",
118 => x"0e3c",
119 => x"0cd6",
120 => x"0b6e",
121 => x"0a04",
122 => x"0898",
123 => x"072c",
124 => x"05be",
125 => x"044f",
126 => x"02df",
127 => x"0170",
128 => x"0000",
129 => x"fe90",
130 => x"fd20",
131 => x"fbb1",
132 => x"fa42",
133 => x"f8d4",
134 => x"f767",
135 => x"f5fc",
136 => x"f492",
137 => x"f32a",
138 => x"f1c4",
139 => x"f060",
140 => x"eefe",
141 => x"ed9f",
142 => x"ec43",
143 => x"eaea",
144 => x"e994",
145 => x"e842",
146 => x"e6f3",
147 => x"e5a8",
148 => x"e461",
149 => x"e31f",
150 => x"e1e1",
151 => x"e0a7",
152 => x"df73",
153 => x"de43",
154 => x"dd19",
155 => x"dbf4",
156 => x"dad4",
157 => x"d9bb",
158 => x"d8a7",
159 => x"d799",
160 => x"d692",
161 => x"d591",
162 => x"d496",
163 => x"d3a2",
164 => x"d2b5",
165 => x"d1cf",
166 => x"d0f0",
167 => x"d019",
168 => x"cf48",
169 => x"ce80",
170 => x"cdbe",
171 => x"cd05",
172 => x"cc54",
173 => x"cbaa",
174 => x"cb09",
175 => x"ca6f",
176 => x"c9de",
177 => x"c956",
178 => x"c8d5",
179 => x"c85e",
180 => x"c7ee",
181 => x"c788",
182 => x"c72a",
183 => x"c6d5",
184 => x"c689",
185 => x"c645",
186 => x"c60b",
187 => x"c5d9",
188 => x"c5b1",
189 => x"c591",
190 => x"c57b",
191 => x"c56d",
192 => x"c569",
193 => x"c56d",
194 => x"c57b",
195 => x"c591",
196 => x"c5b1",
197 => x"c5d9",
198 => x"c60b",
199 => x"c645",
200 => x"c689",
201 => x"c6d5",
202 => x"c72a",
203 => x"c788",
204 => x"c7ee",
205 => x"c85e",
206 => x"c8d5",
207 => x"c956",
208 => x"c9de",
209 => x"ca6f",
210 => x"cb09",
211 => x"cbaa",
212 => x"cc54",
213 => x"cd05",
214 => x"cdbf",
215 => x"ce80",
216 => x"cf49",
217 => x"d019",
218 => x"d0f0",
219 => x"d1cf",
220 => x"d2b5",
221 => x"d3a2",
222 => x"d496",
223 => x"d591",
224 => x"d692",
225 => x"d79a",
226 => x"d8a7",
227 => x"d9bb",
228 => x"dad5",
229 => x"dbf4",
230 => x"dd19",
231 => x"de44",
232 => x"df73",
233 => x"e0a8",
234 => x"e1e1",
235 => x"e31f",
236 => x"e462",
237 => x"e5a9",
238 => x"e6f3",
239 => x"e842",
240 => x"e994",
241 => x"eaea",
242 => x"ec43",
243 => x"ed9f",
244 => x"eefe",
245 => x"f060",
246 => x"f1c4",
247 => x"f32a",
248 => x"f492",
249 => x"f5fc",
250 => x"f768",
251 => x"f8d5",
252 => x"fa42",
253 => x"fbb1",
254 => x"fd21",
255 => x"fe91",
others => x"0000"
);

begin

mem_busy <= mem_readEnable; -- we're done on the cycle after we serve the read request

process (clk, areset)
begin
    if areset = '1' then
    elsif (clk'event and clk = '1') then
        if (mem_writeEnable = '1') then
            ram(to_integer(unsigned(mem_addr(maxAddrBit-1 downto 0)))) := mem_write;
        end if;
        if (mem_readEnable = '1') then
            mem_read <= ram(to_integer(unsigned(mem_addr(maxAddrBit-1 downto 0))));
        end if;
    end if;
end process;

end dram_arch;
